
module PC(
	input  [31:0] NXT_PC,
	input  		  clk,rst,
	output reg [31:0] PC 
);
	
	always @(posedge clk , negedge rst)
	begin
	if(!rst) 
		PC <= 32'h0000_0000 ;
	else
		PC <= NXT_PC ;
	end
	
endmodule 