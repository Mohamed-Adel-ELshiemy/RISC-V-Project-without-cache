library verilog;
use verilog.vl_types.all;
entity Single_Cycle_Top_Tb is
end Single_Cycle_Top_Tb;
